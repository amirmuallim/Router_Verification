class router_vseqs extends uvm_sequence #(uvm_sequence_item);

	`uvm_object_utils(router_vseqs)

	function new(string name = "router_vseqs");
		super.new;
	endfunction : new

endclass : router_vseqs
